`timescale 1ns / 1ps

module ASIC_backup (
  input      nReset,
  input      Clock,
  input      Mode,
  input      Go,
  input      Enable_f,
  input      Sel_f,
  input      S1,
  input      S2,
  input      [5:0] In,
  output     [5:0] DOut1,
  output     [5:0] DOut2,
  output     [5:0] DOut3,
  output     [5:0] DOut4,
  output     [5:0] DOut5,
  output     [5:0] TOut,
  output reg Dclk
);

parameter N1 = 100;
parameter N2 = 6;
parameter N3 = 84;
parameter N4 = 76;
parameter FL = 40;
parameter N = 4;
parameter M = 5;
parameter DCmax = 100;

logic Inkeep;
logic Inshift;
logic Outkeep;
logic Outshift;
logic SelCLK;
logic Start;
logic Sclk;
logic [N2-1:0][N1-1:0] InData;
logic [N3-1:0] Tdata_in;
logic [N4-1:0] Tdata_out;

logic [FL-1:0] b1_ideal;
logic signed [2:0][N-1:0] but1; 
logic signed [FL+2:0][N-1:0] bua2; 
logic signed [FL-1:0][N-1:0] bua3; 
logic signed [2:0][N-1:0] blt1; 
logic signed [FL+2:0][N-1:0] bla2; 
logic Ready1;
logic Valid_Data1;
logic Ready2;
logic Valid_Data2;
logic Ready3;
logic Valid_Data3;
logic Ready4;
logic Valid_Data4;
logic Ready5;
logic Valid_Data5;

reg [N2-1:0][N1-1:0] BusData;

always @ (posedge Clock, negedge nReset) begin
  if (!nReset) begin
    BusData <= 'b0;
  end
  else begin
    if (!Inkeep)
        BusData <= BusData;
    else
		BusData <= InData;
  end
end

assign Tdata_in = InData[0][N3-1:0];

genvar i, j;

for (i=0;i<3;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign but1[i][j] = BusData[0][N*(i)+j];
	end
end

for (i=0;i<22;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bua2[i][j] = BusData[0][N*(i+3)+j];
	end
end

for (i=0;i<FL+3-22;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bua2[i+22][j] = BusData[1][N*(i)+j];
	end
end

for (i=0;i<25-(FL+3-22);i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bua3[i][j] = BusData[1][N*(i+FL+3-22)+j];
	end
end

for (i=0;i<25;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bua3[i+25-(FL+3-22)][j] = BusData[2][N*(i)+j];
	end
end

for (i=0;i<FL+FL-69;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bua3[i+69-FL][j] = BusData[3][N*(i)+j];
	end
end

for (i=0;i<3;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign blt1[i][j] = BusData[3][N*(i+FL+FL-69)+j];
	end
end

for (i=0;i<25-(FL+FL-69+3);i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bla2[i][j] = BusData[3][N*(i+FL+FL-69+3)+j];
	end
end

for (i=0;i<25;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bla2[i+25-(FL+FL-69+3)][j] = BusData[4][N*(i)+j];
	end
end

//25-(FL+FL-69+3)+25=116-FL-FL
//FL+3-(116-FL-FL)=3*FL-113
for (i=0;i<3*FL-113;i++)
begin
	for (j=0;j<4;j++)
	begin
	assign bla2[i+116-FL-FL][j] = BusData[5][N*(i)+j];
	end
end

for (j=0;j<FL;j++)
begin
assign b1_ideal[j] = BusData[5][N*(3*FL-113)+j];
end


SysControl #(.N1(N1), .N2(N2))
SysControl1 (
  .nReset(nReset),
  .Clock(Clock),
  .Mode(Mode),
  .Go(Go),
  .Enable_f(Enable_f),
  .Sel_f(Sel_f),
  .Start(Start),
  .Inkeep(Inkeep),
  .Inshift(Inshift),
  .Outkeep(Outkeep),
  .Outshift(Outshift),
  .SelCLK(SelCLK)
);

divider divider1 (.nReset(nReset), .Clock(Clock), .Sel(SelCLK), .ClockOut(Dclk));

assign Sclk = Enable_f ? Dclk : Clock;

InShiftReg #(.N1(N1), .N2(N2))
InShiftReg1 (.nReset(nReset), .Clock(Sclk), .SelShift(Inshift), .SelKeep(Inkeep), .In(In), .Out(InData));

OutShiftReg #(.N1(N4), .N2(N2))
OutShiftReg1 (.nReset(nReset), .Clock(Clock), .SelShift(Outshift), .SelKeep(Outkeep), .In(Tdata_out), .Out(TOut));

Tmodel #(.N(N), .M(M), .N1(N3), .N2(N4))
tmodel (
 .IN(Tdata_in),
 .S1(S1),
 .S2(S2),
 .Clock(Clock),
 .nReset(nReset),
 .OUT(Tdata_out)
 );

FPTD #(.FL(FL), .DCmax(DCmax), .N(N), .M(M)) 
FPTD1            (.Clock(Clock), 
                  .nReset(nReset), 
                  .Start(Start), 
                  .b1_ideal(b1_ideal),
                  .but1(but1), 
                  .bua2(bua2), 
                  .bua3(bua3), 
                  .blt1(blt1), 
                  .bla2(bla2), 
                  .Ready(Ready1),
                  .Valid_Data(Valid_Data1),
                  .Errors(DOut1));
				  
FPTD #(.FL(FL), .DCmax(DCmax), .N(N), .M(M)) 
FPTD2            (.Clock(Clock), 
                  .nReset(nReset), 
                  .Start(Start), 
                  .b1_ideal(b1_ideal),
                  .but1(but1), 
                  .bua2(bua2), 
                  .bua3(bua3), 
                  .blt1(blt1), 
                  .bla2(bla2), 
                  .Ready(Ready2),
                  .Valid_Data(Valid_Data2),
                  .Errors(DOut2));

				  
FPTD #(.FL(FL), .DCmax(DCmax), .N(N), .M(M)) 
FPTD3            (.Clock(Clock), 
                  .nReset(nReset), 
                  .Start(Start), 
                  .b1_ideal(b1_ideal),
                  .but1(but1), 
                  .bua2(bua2), 
                  .bua3(bua3), 
                  .blt1(blt1), 
                  .bla2(bla2), 
                  .Ready(Ready3),
                  .Valid_Data(Valid_Data3),
                  .Errors(DOut3));				  
				  
FPTD #(.FL(FL), .DCmax(DCmax), .N(N), .M(M)) 
FPTD4            (.Clock(Clock), 
                  .nReset(nReset), 
                  .Start(Start), 
                  .b1_ideal(b1_ideal),
                  .but1(but1), 
                  .bua2(bua2), 
                  .bua3(bua3), 
                  .blt1(blt1), 
                  .bla2(bla2), 
                  .Ready(Ready4),
                  .Valid_Data(Valid_Data4),
                  .Errors(DOut4));				  
				  
FPTD #(.FL(FL), .DCmax(DCmax), .N(N), .M(M)) 
FPTD5            (.Clock(Clock), 
                  .nReset(nReset), 
                  .Start(Start), 
                  .b1_ideal(b1_ideal),
                  .but1(but1), 
                  .bua2(bua2), 
                  .bua3(bua3), 
                  .blt1(blt1), 
                  .bla2(bla2), 
                  .Ready(Ready5),
                  .Valid_Data(Valid_Data5),
                  .Errors(DOut5));
				  
endmodule